module tabla1e1();



endmodule